module bit32Adder( input logic [63:0] operA,operB,output logic [63:0] out);
assign out = operA+operB;
endmodule 