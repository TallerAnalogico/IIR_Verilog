module addUnit(input logic  [31:0] opA,opB,
					output logic [31:0] out);
					
					assign out = opA+opB;
					
endmodule
					