module fixPointMult_tb();

logic [31:0] a_i,b_i,c_o;


fixPointMult DUT(.*);


initial 
	begin
	a_i=32'b00000000000000000000110011001100; //0.05
	b_i=32'b11111111111111111100110011001101; //-0.2
	#1;
	$display("1 result: %b", c_o);
	#1;
	
	a_i=32'b00000000000000000011001100110011;// 0.2
	b_i=32'b11111111111111111100110011001101;//-0.2
	#1;
	$display("2 result: %b", c_o);
	#1;
	
	
	a_i=32'b00000000000001010000000000000000;// 5
	b_i=32'b11111111111111111000000000000000;//-0.5
	#1;
	$display("3 result: %b", c_o);
	#1;
		
	a_i=32'b00000000000001010000000000000000;// 5
	b_i=32'b00000000000000001000000000000000;//0.5
	#1;
	$display("4 result: %b", c_o);
	#1;	

	a_i=32'b11111111111110110000000000000000;// -5
	b_i=32'b11111111111111111011111001011101;// -0.2564
	#1;
	$display("5 result: %b", c_o);
	#1;
	
	
	
	

	end





endmodule