module Top(input logic A,output logic B);
assign B=A ;

endmodule 