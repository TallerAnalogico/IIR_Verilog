  
module xorgate(input logic  signA, signB ,
				output logic result);
				
				assign result = signA^signB;
				
endmodule 